// video_sync_generator.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module video_sync_generator (
		input  wire        video_sync_generator_0_clk_clk,           //       video_sync_generator_0_clk.clk
		input  wire        video_sync_generator_0_clk_reset_reset_n, // video_sync_generator_0_clk_reset.reset_n
		output wire        video_sync_generator_0_in_ready,          //        video_sync_generator_0_in.ready
		input  wire        video_sync_generator_0_in_valid,          //                                 .valid
		input  wire [23:0] video_sync_generator_0_in_data,           //                                 .data
		input  wire        video_sync_generator_0_in_endofpacket,    //                                 .endofpacket
		input  wire        video_sync_generator_0_in_startofpacket,  //                                 .startofpacket
		input  wire        video_sync_generator_0_in_empty,          //                                 .empty
		output wire [23:0] video_sync_generator_0_sync_RGB_OUT,      //      video_sync_generator_0_sync.RGB_OUT
		output wire        video_sync_generator_0_sync_HD,           //                                 .HD
		output wire        video_sync_generator_0_sync_VD,           //                                 .VD
		output wire        video_sync_generator_0_sync_DEN           //                                 .DEN
	);

	altera_avalon_video_sync_generator #(
		.DATA_STREAM_BIT_WIDTH (24),
		.BEATS_PER_PIXEL       (1),
		.NUM_COLUMNS           (1024),
		.NUM_ROWS              (768),
		.H_BLANK_PIXELS        (160),
		.H_FRONT_PORCH_PIXELS  (24),
		.H_SYNC_PULSE_PIXELS   (136),
		.H_SYNC_PULSE_POLARITY (0),
		.V_BLANK_LINES         (29),
		.V_FRONT_PORCH_LINES   (3),
		.V_SYNC_PULSE_LINES    (6),
		.V_SYNC_PULSE_POLARITY (0),
		.TOTAL_HSCAN_PIXELS    (1344),
		.TOTAL_VSCAN_LINES     (806)
	) video_sync_generator_0 (
		.clk     (video_sync_generator_0_clk_clk),           //       clk.clk
		.reset_n (video_sync_generator_0_clk_reset_reset_n), // clk_reset.reset_n
		.ready   (video_sync_generator_0_in_ready),          //        in.ready
		.valid   (video_sync_generator_0_in_valid),          //          .valid
		.data    (video_sync_generator_0_in_data),           //          .data
		.eop     (video_sync_generator_0_in_endofpacket),    //          .endofpacket
		.sop     (video_sync_generator_0_in_startofpacket),  //          .startofpacket
		.empty   (video_sync_generator_0_in_empty),          //          .empty
		.RGB_OUT (video_sync_generator_0_sync_RGB_OUT),      //      sync.export
		.HD      (video_sync_generator_0_sync_HD),           //          .export
		.VD      (video_sync_generator_0_sync_VD),           //          .export
		.DEN     (video_sync_generator_0_sync_DEN)           //          .export
	);

endmodule
